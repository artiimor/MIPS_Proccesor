--------------------------------------------------------------------------------
-- Unidad de control principal del micro. Arq0 2019-2020
--
-- Aitor Melero y Arturo Morcillo 1361
--
--------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity control_unit is
   port (
      -- Entrada = codigo de operacion en la instruccion:
      OpCode  : in  std_logic_vector (5 downto 0); --Cosas que comprobamos (input)
      -- Seniales para el PC
      Branch : out  std_logic; -- 1 = Ejecutandose instruccion branch
      -- Seniales relativas a la memoria
      MemToReg : out  std_logic; -- 1 = Escribir en registro la salida de la mem.
      MemWrite : out  std_logic; -- Escribir la memoria
      MemRead  : out  std_logic; -- Leer la memoria
      -- Seniales para la ALU
      ALUSrc : out  std_logic;                     -- 0 = oper.B es registro, 1 = es valor inm.
      ALUOp  : out  std_logic_vector (2 downto 0); -- Tipo operacion para control de la ALU
      -- Seniales para el GPR
      RegWrite : out  std_logic; -- 1=Escribir registro
      RegDst   : out  std_logic  -- 0=Reg. destino es rt, 1=rd
   );
end control_unit;

architecture rtl of control_unit is

   -- Tipo para los codigos de operacion:
   subtype t_opCode is std_logic_vector (5 downto 0);

   -- Codigos de operacion para las diferentes instrucciones:
   constant OP_RTYPE  : t_opCode := "000000";
   constant OP_BEQ    : t_opCode := "000100";
   constant OP_SW     : t_opCode := "101011";
   constant OP_LW     : t_opCode := "100011";
   constant OP_LUI    : t_opCode := "001111";
   constant OP_ADDI   : t_opCode := "001000";
   constant OP_SLTI   : t_opCode := "001010";
   constant OP_J      : t_opCode := "000010";

begin
    process(OpCode) begin
        case OpCode is
            when OP_RTYPE =>
                Branch <= '0';
                MemToReg <= '0';
                MemWrite <= '0';
                ALUSrc <= '0';
                ALUOp <= "111"; --Para el caso de las R tenemos el 111
                RegWrite <= '1';
                MemRead <= '0';
                RegDst <= '1'; -- el unico con 1 obligatorio. El resto operan con datos inmediatos
   
           when OP_BEQ =>
               Branch <= '0'; -- Es un salto
               MemToReg <= '0'; -- Da igual porque regwrite es 0
               MemWrite <= '0';
               ALUSrc <= '0';
               ALUOp <= "001"; --Para el beq ponemos 001 que nos realiza directamente una resta
               RegWrite <= '0';
               MemRead <= '0';
               RegDst <= '0'; --da igual porque regwrite es 0
 
           when OP_SW =>
               Branch <= '0';
               MemToReg <= '0'; -- Da igual porque regwrite es 0
               MemWrite <= '1';
               ALUSrc <= '1';
               ALUOp <= "000"; -- Para que la ALU directamtente sume 000
               RegWrite <= '0';
               MemRead <= '0';
               RegDst <= '1'; --da igual porque regwrite es 0

           when OP_LW =>
               Branch <= '0';
               MemToReg <= '1';
               MemWrite <= '0';
               ALUSrc <= '1'; 
               ALUOp <= "000"; -- Para que la ALU directamtente sume 000
               RegWrite <= '1';
               MemRead <= '1';
               RegDst <= '0';

            when OP_ADDI =>
                Branch <= '0';
                MemToReg <= '0'; --da igual
                MemWrite <= '0';
                ALUSrc <= '1'; --operacion con el inmediato
                ALUOp <= "000"; --Para que la alu sume directamente un 000
                RegWrite <= '1';
                MemRead <= '0';
                RegDst <= '0';
            when OP_LUI =>
                Branch <= '0';
                MemToReg <= '0';
                MemWrite <= '0';
                ALUSrc <= '1'; --En la alu queremos el inmediato
                ALUOp <=  "010";--para lui 010
                RegWrite <= '1';
                MemRead <= '0'; --da igual
                RegDst <= '0';

            when OP_SLTI =>
                Branch <= '0';
                MemToReg <= '0'; --da igual
                MemWrite <= '0';
                ALUSrc <= '1'; --operacion con el inmediato
                ALUOp <=  "011";--para slti 011
                RegWrite <= '1';
                MemRead <= '0';
                RegDst <= '0';

            when OP_J =>
                Branch <= '0';
                MemToReg <= '0';
                MemWrite <= '0';
                ALUSrc <= '1';
                ALUOp <= "100";-- para j quiero el 100
                RegWrite <= '0';
                MemRead <= '0';
                RegDst <= '0';

            when others => --Para el nop
                Branch <= '0';
                MemToReg <= '0';
                MemWrite <= '0';
                ALUSrc <= '0';
                ALUOp <= "111";
                RegWrite <= '0';
                MemRead <= '0';
                RegDst <= '0';
        end case;
    end process;
end architecture;